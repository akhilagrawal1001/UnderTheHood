module or(a,b,c);
intput a,b;
output c;
xnor(c,a,b);
endmodule