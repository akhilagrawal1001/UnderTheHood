module or(a,b,c);
intput a,b;
output c;
or(c,a,b);
endmodule